module ativador( RHX00, RHX01, RHX02, RHX03, RHX04, RHX05, RHX06,
				RHX10, RHX11, RHX12, RHX13, RHX14, RHX15, RHX16,
				RHX20, RHX21, RHX22, RHX23, RHX24, RHX25, RHX26,
				RHX30, RHX31, RHX32, RHX33, RHX34, RHX35, RHX36,
				RHX40, RHX41, RHX42, RHX43, RHX44, RHX45, RHX46,
				RHX50, RHX51, RHX52, RHX53, RHX54, RHX55, RHX56,
				RHX60, RHX61, RHX62, RHX63, RHX64, RHX65, RHX66,
				RHX70, RHX71, RHX72, RHX73, RHX74, RHX75, RHX76,
				
				CHX00, CHX01, CHX02, CHX03, CHX04, CHX05, CHX06,
				CHX10, CHX11, CHX12, CHX13, CHX14, CHX15, CHX16,
				CHX20, CHX21, CHX22, CHX23, CHX24, CHX25, CHX26,
				CHX30, CHX31, CHX32, CHX33, CHX34, CHX35, CHX36,
				CHX40, CHX41, CHX42, CHX43, CHX44, CHX45, CHX46,
				CHX50, CHX51, CHX52, CHX53, CHX54, CHX55, CHX56,
				CHX60, CHX61, CHX62, CHX63, CHX64, CHX65, CHX66,
				CHX70, CHX71, CHX72, CHX73, CHX74, CHX75, CHX76,
				seletor, clock,
				SHX00, SHX01, SHX02, SHX03, SHX04, SHX05, SHX06,
				SHX10, SHX11, SHX12, SHX13, SHX14, SHX15, SHX16,
				SHX20, SHX21, SHX22, SHX23, SHX24, SHX25, SHX26,
				SHX30, SHX31, SHX32, SHX33, SHX34, SHX35, SHX36,
				SHX40, SHX41, SHX42, SHX43, SHX44, SHX45, SHX46,
				SHX50, SHX51, SHX52, SHX53, SHX54, SHX55, SHX56,
				SHX60, SHX61, SHX62, SHX63, SHX64, SHX65, SHX66,
				SHX70, SHX71, SHX72, SHX73, SHX74, SHX75, SHX76);
input seletor, clock;
input 	RHX00, RHX01, RHX02, RHX03, RHX04, RHX05, RHX06,
		RHX10, RHX11, RHX12, RHX13, RHX14, RHX15, RHX16,
		RHX20, RHX21, RHX22, RHX23, RHX24, RHX25, RHX26,
		RHX30, RHX31, RHX32, RHX33, RHX34, RHX35, RHX36,
		RHX40, RHX41, RHX42, RHX43, RHX44, RHX45, RHX46,
		RHX50, RHX51, RHX52, RHX53, RHX54, RHX55, RHX56,
		RHX60, RHX61, RHX62, RHX63, RHX64, RHX65, RHX66,
		RHX70, RHX71, RHX72, RHX73, RHX74, RHX75, RHX76,		
		CHX00, CHX01, CHX02, CHX03, CHX04, CHX05, CHX06,
		CHX10, CHX11, CHX12, CHX13, CHX14, CHX15, CHX16,
		CHX20, CHX21, CHX22, CHX23, CHX24, CHX25, CHX26,
		CHX30, CHX31, CHX32, CHX33, CHX34, CHX35, CHX36,
		CHX40, CHX41, CHX42, CHX43, CHX44, CHX45, CHX46,
		CHX50, CHX51, CHX52, CHX53, CHX54, CHX55, CHX56,
		CHX60, CHX61, CHX62, CHX63, CHX64, CHX65, CHX66,
		CHX70, CHX71, CHX72, CHX73, CHX74, CHX75, CHX76;
	
output reg 	SHX00, SHX01, SHX02, SHX03, SHX04, SHX05, SHX06,
			SHX10, SHX11, SHX12, SHX13, SHX14, SHX15, SHX16,
			SHX20, SHX21, SHX22, SHX23, SHX24, SHX25, SHX26,
			SHX30, SHX31, SHX32, SHX33, SHX34, SHX35, SHX36,
			SHX40, SHX41, SHX42, SHX43, SHX44, SHX45, SHX46,
			SHX50, SHX51, SHX52, SHX53, SHX54, SHX55, SHX56,
			SHX60, SHX61, SHX62, SHX63, SHX64, SHX65, SHX66,
			SHX70, SHX71, SHX72, SHX73, SHX74, SHX75, SHX76;

always @(posedge clock) begin
	case(seletor)
		1 : begin 
				SHX00 = CHX00; SHX01 = CHX01; SHX02 = CHX02; SHX03 = CHX03; SHX04 = CHX04; SHX05 = CHX05; SHX06 = CHX06;
				SHX10 = CHX10; SHX11 = CHX11; SHX12 = CHX12; SHX13 = CHX13; SHX14 = CHX14; SHX15 = CHX15; SHX16 = CHX16;
				SHX20 = CHX20; SHX21 = CHX21; SHX22 = CHX22; SHX23 = CHX23; SHX24 = CHX24; SHX25 = CHX25; SHX26 = CHX26;
				SHX30 = CHX30; SHX31 = CHX31; SHX32 = CHX32; SHX33 = CHX33; SHX34 = CHX34; SHX35 = CHX35; SHX36 = CHX36;
				SHX40 = CHX40; SHX41 = CHX41; SHX42 = CHX42; SHX43 = CHX43; SHX44 = CHX44; SHX45 = CHX45; SHX46 = CHX46;
				SHX50 = CHX50; SHX51 = CHX51; SHX52 = CHX52; SHX53 = CHX53; SHX54 = CHX54; SHX55 = CHX55; SHX56 = CHX56;
				SHX60 = CHX60; SHX61 = CHX61; SHX62 = CHX62; SHX63 = CHX63; SHX64 = CHX64; SHX65 = CHX65; SHX66 = CHX66;
				SHX70 = CHX70; SHX71 = CHX71; SHX72 = CHX72; SHX73 = CHX73; SHX74 = CHX74; SHX75 = CHX75; SHX76 = CHX76;
			end
		0 : begin 
				SHX00 = RHX00; SHX01 = RHX01; SHX02 = RHX02; SHX03 = RHX03; SHX04 = RHX04; SHX05 = RHX05; SHX06 = RHX06;
				SHX10 = RHX10; SHX11 = RHX11; SHX12 = RHX12; SHX13 = RHX13; SHX14 = RHX14; SHX15 = RHX15; SHX16 = RHX16;
				SHX20 = RHX20; SHX21 = RHX21; SHX22 = RHX22; SHX23 = RHX23; SHX24 = RHX24; SHX25 = RHX25; SHX26 = RHX26;
				SHX30 = RHX30; SHX31 = RHX31; SHX32 = RHX32; SHX33 = RHX33; SHX34 = RHX34; SHX35 = RHX35; SHX36 = RHX36;
				SHX40 = RHX40; SHX41 = RHX41; SHX42 = RHX42; SHX43 = RHX43; SHX44 = RHX44; SHX45 = RHX45; SHX46 = RHX46;
				SHX50 = RHX50; SHX51 = RHX51; SHX52 = RHX52; SHX53 = RHX53; SHX54 = RHX54; SHX55 = RHX55; SHX56 = RHX56;
				SHX60 = RHX60; SHX61 = RHX61; SHX62 = RHX62; SHX63 = RHX63; SHX64 = RHX64; SHX65 = RHX65; SHX66 = RHX66;
				SHX70 = RHX70; SHX71 = RHX71; SHX72 = RHX72; SHX73 = RHX73; SHX74 = RHX74; SHX75 = RHX75; SHX76 = RHX76;
			end
	endcase
end
endmodule
